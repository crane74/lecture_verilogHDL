/* 1 bit and */

module and (input a, b, output s );

  assign s = a & b  ;  // adder.vの+を&に変えただけ

endmodule



