/* 1 bit adder */

module adder (input a, b, output s );

  assign s = a + b  ;  // add a b

endmodule



